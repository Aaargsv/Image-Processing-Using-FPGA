module image_proc_top_design
	(
		input  logic 			i_clk,
		input  logic 			i_reset_n,
		input  logic 			i_pclk,
		input  logic [7 : 0]	i_data,
		input  logic 			i_hsync,
		input  logic			i_vsync,
		input  logic 			i_red_screen,

		input  logic			i_change_kernel,
		input  logic 			i_select_mode,
		input  logic			i_threshold,

		output logic 			o_device_working,
		output logic 			o_xclk,
		output logic			o_siod,
		output logic			o_sioc,

		output logic 		 	o_vga_hsync,
		output logic 		 	o_vga_vsync,
		output logic [7 : 0]	o_vga_r,
		output logic [7 : 0]	o_vga_g,
		output logic [7 : 0]	o_vga_b,
		output logic 			o_dac_nblank,
		output logic  			o_dac_clk,
		output logic 			o_dac_nsync,
		output logic 			o_camera_reset,
		output logic			o_camera_pwdn

	);


	localparam FREQ_GLOBAL		   		= 50_000_000;
	localparam FREQ_CAM		       		= 25_000_000;
	localparam FREQ_SCCB				= 100000;

	localparam KERNEL 			  	    = 3;
	localparam KERNEL_NUM_ELEMENTS 		= KERNEL * KERNEL;
	localparam COLOR_CHANNEL	   		= 8;
	localparam WIDTH_IMAGE		   		= 640;
	localparam HEIGHT_IMAGE				= 480;
	localparam DATA_KERNEL_WIDTH		= COLOR_CHANNEL + 1;

	localparam MEM_DEPTH = 262144;

	logic signed   [DATA_KERNEL_WIDTH   - 1 : 0]   	w_kernel   			  [1 : 0][KERNEL_NUM_ELEMENTS  - 1 : 0];
	logic signed   [DATA_KERNEL_WIDTH   - 1 : 0]   	w_kernel_from_mem            [KERNEL_NUM_ELEMENTS  - 1 : 0];

	logic		      [15 : 0]								   w_pixel_data_16;
	logic		      [18 : 0]								   wr_address;


	logic			w_clk_50mhz;
	logic 			w_clk_25mhz;
	logic 			w_config_done;
	logic 			w_config_start;
	logic 			w_device_work_start;

	logic 			w_pixel_ready;
	logic 			w_pixel_data_valid;

	logic			[15 : 0]	wr_ram_data;
	logic			[18 : 0]	rd_address_ram_to_vga;
	logic 			[2  : 0]	w_kernel_address;

	logic			w_we_memory;

	logic w_sioc;
	logic w_siod;
	assign o_sioc 			= w_sioc ? 1'b1 : 1'b0;
	assign o_siod 			= w_siod ? 1'b1 : 1'b0;

	assign dac_nsync      = 1'bz;
	assign o_camera_pwdn  = 1'b0;

	assign o_xclk 			= w_clk_25mhz;
	assign w_clk_50mhz 		= i_clk;
	assign o_device_working = w_device_work_start;
	assign o_camera_reset 	= i_reset_n;


	address_kernel_counter address_kernel_counter_inst
	(
		.i_clk		(w_clk_50mhz),
		.i_reset_n	(i_reset_n),
		.i_button	(i_change_kernel),

		.o_address	(w_kernel_address)

	);

	kernel_mem
	#(
		.KERNEL_NUM_ELEMENTS (KERNEL_NUM_ELEMENTS),
		.DATA_KERNEL_WIDTH   (DATA_KERNEL_WIDTH)
	)
		kernel_mem_inst
	(
			.i_clk 				(i_clk),
			.i_kernel_address	(i_kernel_address),
			.o_kernel			(w_kernel_from_mem)
	);


	logic w_select_mode;
	logic w_threshold;


	assign w_threshold   = ~i_threshold;
	assign w_select_mode = ~i_select_mode;

	/*selection_mode selection_mode_inst
	(
		.i_clk			(i_clk),
		.i_reset_n		(i_reset_n),
		.i_select_mode	(i_select_mode),

		.o_select_mode	(w_select_mode),
		.o_threshold	(w_threshold)
	);*/

	always_comb
		begin
			if (w_select_mode)
				w_kernel[0] = '{ 	-1,  0, 1,
									-2,  0, 2,
									-1,  0, 1 };
			else
				w_kernel[0] = w_kernel_from_mem;
		end


	assign w_kernel[1] =  '{ -1,  -2, -1,
							  0,   0,  0,
							  1,   2,  1 };


	clock_divider
	#(
		.FREQ_1	(FREQ_GLOBAL),
		.FREQ_2	(FREQ_CAM)
	)
	clock_divider_inst
	(
		 .i_clk		(w_clk_50mhz),
		 .i_reset_n (i_reset_n),
		 .o_clk		(w_clk_25mhz)
	);

	main_control main_control_inst
	(
		 .i_clk					(w_clk_25mhz),
		 .i_reset_n				(i_reset_n),
		 .i_config_done			(w_config_done),
		 .o_config_start		(w_config_start),
		 .o_device_work_start	(w_device_work_start)
	);

	camera_configuration
	#(
	.CLK_FREQUENCY		(FREQ_CAM),
	.SCCB_FREQUENCY 	(FREQ_SCCB)
	)
	camera_configuration_inst
	(
		.i_clk			(w_clk_25mhz),
		.i_reset_n		(i_reset_n),
		.i_config_start	(w_config_start),

		.o_config_done	(w_config_done),
		.o_sioc			(w_sioc),
		.o_siod			(w_siod)
	);



	pixel_capture #(.MAX_ADDRESS(MEM_DEPTH - 1))
	pixel_capture_inst
	(
		.i_clk					(w_clk_50mhz),
		.i_pclk					(i_pclk),
		.i_reset_n				(i_reset_n),
		.i_data					(i_data),
		.i_hsync				(i_hsync),
		.i_vsync				(i_vsync),
		.i_device_work_start	(w_device_work_start),
		.o_pixel_data			(w_pixel_data_16),
		.o_pixel_ready			(w_pixel_ready),

		.o_we_memory			(w_we_memory),
		.o_vsync                (),
		.o_fake_output			(),
		.o_wr_address           ()
	);


	logic [2 : 0][COLOR_CHANNEL - 1 : 0] 					w_data_from_wb [1 : 0];
	logic [KERNEL - 1 : 0][2 : 0][COLOR_CHANNEL - 1 : 0] 	w_pixel_area_data 		   [KERNEL - 1 : 0];
	logic 													w_pixel_data_valid_wb;

	logic [2 : 0][COLOR_CHANNEL - 1 : 0] 					w_data_from_mux;
	logic 								 					w_data_ready_from_mux;
	logic [2 : 0][COLOR_CHANNEL - 1 : 0] 					w_data_to_ram;
	logic 								 					w_wr_enable;
	logic [COLOR_CHANNEL - 1 : 0]		   					w_convolution_value		   [1 : 0][2 : 0];
	logic [2 : 0][COLOR_CHANNEL - 1 : 0]					w_magnitude_value;
	logic													w_magnitude_ready;

	window_buffer
	#(
		.COLOR_CHANNEL	(COLOR_CHANNEL),
		.KERNEL		  	(KERNEL),
		.WIDTH_IMAGE  	(WIDTH_IMAGE),
		.HEIGHT_IMAGE	(HEIGHT_IMAGE)

	) window_buffer_inst
	  (
		.i_clk						(w_clk_50mhz),
		.i_reset_n					(i_reset_n),
		.i_pixel_data				({	w_pixel_data_16[15 : 11], w_pixel_data_16[15 : 13],
									    w_pixel_data_16[10 : 5],  w_pixel_data_16[10 : 9],
			                            w_pixel_data_16[4  : 0],  w_pixel_data_16[4  : 2]
									}),

		.i_pixel_ready			(w_pixel_ready),
		.o_pixel_area_data		(w_pixel_area_data),
		.o_pixel_data_valid		(w_pixel_data_valid_wb)
	);



	convolution_set
	#(
		.KERNEL					(KERNEL),
		.KERNEL_NUM_ELEMENTS	(KERNEL_NUM_ELEMENTS),
		.COLOR_CHANNEL			(COLOR_CHANNEL),
		.DATA_KERNEL_WIDTH		(DATA_KERNEL_WIDTH)
	)
	convolution_set_inst_0
	(
		.i_kernel   			(w_kernel[0]),
		.i_pixel_area_data 		(w_pixel_area_data),
		.o_convolution_value	(w_convolution_value[0])
	);

	convolution_set
	#(
		.KERNEL					(KERNEL),
		.KERNEL_NUM_ELEMENTS	(KERNEL_NUM_ELEMENTS),
		.COLOR_CHANNEL			(COLOR_CHANNEL),
		.DATA_KERNEL_WIDTH		(DATA_KERNEL_WIDTH)
	)
	convolution_set_inst_1
	(
		.i_kernel   			(w_kernel[1]),
		.i_pixel_area_data 		(w_pixel_area_data),
		.o_convolution_value	(w_convolution_value[1])

	);

	magnitude
	#(
		.COLOR_CHANNEL (COLOR_CHANNEL)
	)
	magnitude_inst
	(
		.i_clk					(i_clk),
		.i_reset_n				(i_reset_n),
		.i_data_ready			(w_pixel_data_valid_wb),
		.i_convolution_value	(w_convolution_value),

		.o_data_ready			(w_magnitude_ready),
		.o_magnitude_value		(w_magnitude_value)
	);

	 mux#(.COLOR_CHANNEL(COLOR_CHANNEL))
	 mux_inst
	(
		.i_select_mode						(w_select_mode),

		.i_single_filter_convolution_value 	(w_convolution_value[0]),
		.i_magnitude_value					(w_magnitude_value),

		.i_signle_filter_data_ready			(w_pixel_data_valid_wb),
		.i_magnitude_data_ready				(w_magnitude_ready),

		.o_data								(w_data_from_mux),
		.o_data_ready						(w_data_ready_from_mux)
	);


	logic [2 : 0][COLOR_CHANNEL - 1 : 0]    w_post_proc_data;
	logic									w_post_proc_ready;

	post_proc #(.COLOR_CHANNEL(COLOR_CHANNEL)) post_proc_inst
	(
		.i_clk				(i_clk),
		.i_reset_n			(i_reset_n),

		.i_data_ready		(w_data_ready_from_mux),
		.i_data				(w_data_from_mux),
		.i_kernel_address	(w_kernel_address),
		.i_select_mode		(w_select_mode),
		.i_threshold		(w_threshold),

		.o_data_ready		(w_post_proc_ready),
		.o_data				(w_post_proc_data)

	);


	writer
	#(
		.MAX_ADDRESS	(MEM_DEPTH - 1),
		.COLOR_CHANNEL	(COLOR_CHANNEL),
		.WIDTH_IMAGE	(WIDTH_IMAGE),
		.HEIGHT_IMAGE	(HEIGHT_IMAGE)
	)
	writer_inst
	(
		.i_clk			(w_clk_50mhz),
		.i_data_ready	(w_post_proc_ready),
		.i_reset_n		(i_reset_n),
		.i_data			(w_post_proc_data),

		.o_wr_enable    (w_wr_enable),
		.o_data			(w_data_to_ram),
		.o_wr_address	(wr_address)
	);


	RAM_16 #( .DEPTH(MEM_DEPTH))
	RAM_16_inst
	(
		 .i_clk					(w_clk_50mhz),
		 .i_write_enable 		(w_wr_enable),
		 .i_write_address		(wr_address			    [$clog2(MEM_DEPTH) - 1 : 0]),
		 .i_read_address		(rd_address_ram_to_vga	[$clog2(MEM_DEPTH) - 1 : 0]),
		 .i_write_value 
		 (
			{	w_data_to_ram[2][7 : 3],
				w_data_to_ram[1][7 : 2],
				w_data_to_ram[0][7 : 3]
			}
		 ),
		 .o_read_value			(wr_ram_data)
	);

	
	VGA VGA_inst
		(
			.i_clk				(w_clk_25mhz),
			.i_data				(wr_ram_data),
			.i_reset_n			(i_reset_n),

			.i_red_screen		(i_red_screen),

			.o_pixel_counter	(rd_address_ram_to_vga),
			.o_hsync				(o_vga_hsync),
			.o_vsync				(o_vga_vsync),
			.o_R					(o_vga_r),
			.o_G					(o_vga_g),
			.o_B					(o_vga_b),

			.o_clk				(o_dac_clk),
			.o_nsync			(o_dac_nsync),
			.o_nblank			(o_dac_nblank)
		);

endmodule : image_proc_top_design
