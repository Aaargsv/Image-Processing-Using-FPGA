module mux
    #(
        parameter COLOR_CHANNEL
    )
    (
        input   logic i_select_mode,

        input   logic [COLOR_CHANNEL - 1 : 0]	        i_single_filter_convolution_value [2 : 0],
        input   logic [2 : 0][COLOR_CHANNEL - 1 : 0]    i_magnitude_value,

        input   logic                                   i_signle_filter_data_ready,
        input   logic                                   i_magnitude_data_ready,

        output  logic [2 : 0][COLOR_CHANNEL - 1 : 0]    o_data,
        output  logic                                   o_data_ready
    );

    assign o_data       = (i_select_mode) ? (i_magnitude_value)         : {i_single_filter_convolution_value[2], 
																									i_single_filter_convolution_value[1],
																									i_single_filter_convolution_value[0]};
																									
    assign o_data_ready = (i_select_mode) ? (i_magnitude_data_ready)    : i_signle_filter_data_ready;


endmodule : mux
